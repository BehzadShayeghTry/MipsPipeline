module Adder(input [4:0] in, pluser, output out);
    assign out = in + pluser;
endmodule