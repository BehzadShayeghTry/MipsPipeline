module Adder(input [4:0] in, pluser, output [4:0] out);
    assign out = in + pluser;
endmodule